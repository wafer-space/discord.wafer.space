magic
tech gf180mcuD
magscale 1 10
timestamp 1764882048
<< nwell >>
rect -86 354 4230 870
<< pwell >>
rect -86 -86 4230 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 583 68 639 268
rect 887 68 943 268
rect 1258 68 1314 268
rect 1374 68 1430 268
rect 1516 68 1572 268
rect 1738 68 1794 268
rect 1956 68 2012 268
rect 2204 68 2260 268
rect 2391 68 2447 268
rect 2895 68 2951 268
rect 3062 68 3118 268
rect 3270 68 3326 268
rect 3456 68 3512 268
rect 3777 68 3833 268
rect 3937 68 3993 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 588 440 645 716
rect 777 440 833 716
rect 1061 440 1118 716
rect 1356 440 1412 716
rect 1516 440 1572 716
rect 1807 440 1863 716
rect 2009 440 2065 716
rect 2324 440 2380 716
rect 2509 440 2565 716
rect 2895 440 2951 716
rect 3082 440 3138 716
rect 3270 440 3326 716
rect 3456 440 3512 716
rect 3777 440 3833 716
rect 3937 440 3993 716
<< ndiff >>
rect 28 255 116 268
rect 28 209 41 255
rect 87 209 116 255
rect 28 68 116 209
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 255 429 268
rect 332 209 361 255
rect 407 209 429 255
rect 332 68 429 209
rect 485 127 583 268
rect 485 81 498 127
rect 544 81 583 127
rect 485 68 583 81
rect 639 255 887 268
rect 639 209 682 255
rect 728 209 887 255
rect 639 68 887 209
rect 943 255 1258 268
rect 943 209 986 255
rect 1032 209 1258 255
rect 943 68 1258 209
rect 1314 68 1374 268
rect 1430 68 1516 268
rect 1572 127 1738 268
rect 1572 81 1651 127
rect 1697 81 1738 127
rect 1572 68 1738 81
rect 1794 68 1956 268
rect 2012 255 2204 268
rect 2012 209 2098 255
rect 2144 209 2204 255
rect 2012 68 2204 209
rect 2260 255 2391 268
rect 2260 209 2316 255
rect 2362 209 2391 255
rect 2260 68 2391 209
rect 2447 255 2693 268
rect 2447 209 2634 255
rect 2680 209 2693 255
rect 2447 68 2693 209
rect 2773 255 2895 268
rect 2773 209 2809 255
rect 2855 209 2895 255
rect 2773 68 2895 209
rect 2951 68 3062 268
rect 3118 127 3270 268
rect 3118 81 3195 127
rect 3241 81 3270 127
rect 3118 68 3270 81
rect 3326 68 3456 268
rect 3512 255 3613 268
rect 3512 152 3554 255
rect 3600 152 3613 255
rect 3512 68 3613 152
rect 3689 255 3777 268
rect 3689 81 3702 255
rect 3748 81 3777 255
rect 3689 68 3777 81
rect 3833 255 3937 268
rect 3833 117 3862 255
rect 3908 117 3937 255
rect 3833 68 3937 117
rect 3993 255 4116 268
rect 3993 81 4022 255
rect 4068 81 4116 255
rect 3993 68 4116 81
<< pdiff >>
rect 28 587 116 716
rect 28 541 41 587
rect 87 541 116 587
rect 28 440 116 541
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 499 429 716
rect 332 453 361 499
rect 407 453 429 499
rect 332 440 429 453
rect 485 703 588 716
rect 485 657 498 703
rect 544 657 588 703
rect 485 440 588 657
rect 645 574 777 716
rect 645 468 693 574
rect 739 468 777 574
rect 645 440 777 468
rect 833 569 1061 716
rect 833 453 986 569
rect 1032 453 1061 569
rect 833 440 1061 453
rect 1118 622 1356 716
rect 1118 576 1182 622
rect 1228 576 1356 622
rect 1118 440 1356 576
rect 1412 703 1516 716
rect 1412 657 1441 703
rect 1487 657 1516 703
rect 1412 440 1516 657
rect 1572 625 1663 716
rect 1572 579 1601 625
rect 1647 579 1663 625
rect 1572 440 1663 579
rect 1719 622 1807 716
rect 1719 576 1732 622
rect 1778 576 1807 622
rect 1719 440 1807 576
rect 1863 703 2009 716
rect 1863 657 1909 703
rect 1955 657 2009 703
rect 1863 440 2009 657
rect 2065 499 2324 716
rect 2065 453 2109 499
rect 2155 453 2324 499
rect 2065 440 2324 453
rect 2380 666 2509 716
rect 2380 460 2431 666
rect 2477 460 2509 666
rect 2380 440 2509 460
rect 2565 501 2688 716
rect 2565 455 2611 501
rect 2657 455 2688 501
rect 2565 440 2688 455
rect 2787 703 2895 716
rect 2787 653 2817 703
rect 2863 653 2895 703
rect 2787 440 2895 653
rect 2951 572 3082 716
rect 2951 463 3001 572
rect 3047 463 3082 572
rect 2951 440 3082 463
rect 3138 703 3270 716
rect 3138 656 3186 703
rect 3232 656 3270 703
rect 3138 440 3270 656
rect 3326 573 3456 716
rect 3326 453 3370 573
rect 3416 453 3456 573
rect 3326 440 3456 453
rect 3512 703 3631 716
rect 3512 453 3572 703
rect 3618 453 3631 703
rect 3512 440 3631 453
rect 3689 703 3777 716
rect 3689 453 3702 703
rect 3748 453 3777 703
rect 3689 440 3777 453
rect 3833 667 3937 716
rect 3833 453 3862 667
rect 3908 453 3937 667
rect 3833 440 3937 453
rect 3993 703 4116 716
rect 3993 453 4022 703
rect 4068 453 4116 703
rect 3993 440 4116 453
<< ndiffc >>
rect 41 209 87 255
rect 201 81 247 127
rect 361 209 407 255
rect 498 81 544 127
rect 682 209 728 255
rect 986 209 1032 255
rect 1651 81 1697 127
rect 2098 209 2144 255
rect 2316 209 2362 255
rect 2634 209 2680 255
rect 2809 209 2855 255
rect 3195 81 3241 127
rect 3554 152 3600 255
rect 3702 81 3748 255
rect 3862 117 3908 255
rect 4022 81 4068 255
<< pdiffc >>
rect 41 541 87 587
rect 201 657 247 703
rect 361 453 407 499
rect 498 657 544 703
rect 693 468 739 574
rect 986 453 1032 569
rect 1182 576 1228 622
rect 1441 657 1487 703
rect 1601 579 1647 625
rect 1732 576 1778 622
rect 1909 657 1955 703
rect 2109 453 2155 499
rect 2431 460 2477 666
rect 2611 455 2657 501
rect 2817 653 2863 703
rect 3001 463 3047 572
rect 3186 656 3232 703
rect 3370 453 3416 573
rect 3572 453 3618 703
rect 3702 453 3748 703
rect 3862 453 3908 667
rect 4022 453 4068 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 588 716 645 760
rect 777 716 833 760
rect 1061 716 1118 760
rect 1356 716 1412 760
rect 1516 716 1572 760
rect 1807 716 1863 760
rect 2009 716 2065 760
rect 2324 716 2380 760
rect 2509 716 2565 760
rect 2895 716 2951 760
rect 3082 716 3138 760
rect 3270 716 3326 760
rect 3456 716 3512 760
rect 3777 716 3833 760
rect 3937 716 3993 760
rect 116 394 172 440
rect 100 379 172 394
rect 276 393 332 440
rect 588 398 645 440
rect 777 420 833 440
rect 761 407 833 420
rect 100 333 113 379
rect 159 333 172 379
rect 100 320 172 333
rect 116 268 172 320
rect 222 378 332 393
rect 222 332 235 378
rect 281 332 332 378
rect 222 319 332 332
rect 577 385 649 398
rect 577 339 590 385
rect 636 339 649 385
rect 761 361 774 407
rect 820 361 833 407
rect 1061 398 1118 440
rect 1356 419 1412 440
rect 1061 385 1137 398
rect 1356 395 1430 419
rect 761 348 833 361
rect 881 371 953 384
rect 577 326 649 339
rect 276 268 332 319
rect 583 268 639 326
rect 881 325 894 371
rect 940 325 953 371
rect 1061 339 1078 385
rect 1124 339 1137 385
rect 1374 371 1430 395
rect 1516 371 1572 440
rect 1807 397 1863 440
rect 2009 397 2065 440
rect 2324 397 2380 440
rect 2509 416 2565 440
rect 2509 403 2585 416
rect 1807 393 1877 397
rect 1738 384 1877 393
rect 1061 326 1137 339
rect 1250 347 1322 360
rect 881 312 953 325
rect 887 268 943 312
rect 1250 301 1263 347
rect 1309 301 1322 347
rect 1250 288 1322 301
rect 1374 358 1446 371
rect 1374 312 1387 358
rect 1433 312 1446 358
rect 1374 299 1446 312
rect 1516 358 1589 371
rect 1516 312 1530 358
rect 1576 312 1589 358
rect 1516 299 1589 312
rect 1738 338 1818 384
rect 1864 338 1877 384
rect 2000 384 2076 397
rect 2000 378 2015 384
rect 1738 325 1877 338
rect 1956 338 2015 378
rect 2061 338 2076 384
rect 2324 384 2447 397
rect 1956 325 2076 338
rect 2196 347 2268 360
rect 1258 268 1314 288
rect 1374 268 1430 299
rect 1516 268 1572 299
rect 1738 268 1794 325
rect 1956 268 2012 325
rect 2196 301 2209 347
rect 2255 301 2268 347
rect 2324 338 2339 384
rect 2385 338 2447 384
rect 2509 357 2524 403
rect 2570 357 2585 403
rect 2895 397 2951 440
rect 2509 344 2585 357
rect 2875 384 2951 397
rect 3082 395 3138 440
rect 2324 325 2447 338
rect 2875 338 2888 384
rect 2934 338 2951 384
rect 2875 325 2951 338
rect 2196 288 2268 301
rect 2204 268 2260 288
rect 2391 268 2447 325
rect 2895 268 2951 325
rect 3062 382 3153 395
rect 3062 336 3093 382
rect 3139 336 3153 382
rect 3270 360 3326 440
rect 3062 323 3153 336
rect 3254 347 3326 360
rect 3062 268 3118 323
rect 3254 301 3267 347
rect 3313 301 3326 347
rect 3254 288 3326 301
rect 3270 268 3326 288
rect 3456 420 3512 440
rect 3456 407 3532 420
rect 3456 361 3473 407
rect 3519 361 3532 407
rect 3777 396 3833 440
rect 3937 396 3993 440
rect 3456 348 3532 361
rect 3600 383 3993 396
rect 3456 268 3512 348
rect 3600 337 3624 383
rect 3780 337 3993 383
rect 3600 324 3993 337
rect 3777 268 3833 324
rect 3937 268 3993 324
rect 116 24 172 68
rect 276 24 332 68
rect 583 24 639 68
rect 887 24 943 68
rect 1258 24 1314 68
rect 1374 24 1430 68
rect 1516 24 1572 68
rect 1738 24 1794 68
rect 1956 24 2012 68
rect 2204 24 2260 68
rect 2391 24 2447 68
rect 2895 24 2951 68
rect 3062 24 3118 68
rect 3270 24 3326 68
rect 3456 24 3512 68
rect 3777 24 3833 68
rect 3937 24 3993 68
<< polycontact >>
rect 113 333 159 379
rect 235 332 281 378
rect 590 339 636 385
rect 774 361 820 407
rect 894 325 940 371
rect 1078 339 1124 385
rect 1263 301 1309 347
rect 1387 312 1433 358
rect 1530 312 1576 358
rect 1818 338 1864 384
rect 2015 338 2061 384
rect 2209 301 2255 347
rect 2339 338 2385 384
rect 2524 357 2570 403
rect 2888 338 2934 384
rect 3093 336 3139 382
rect 3267 301 3313 347
rect 3473 361 3519 407
rect 3624 337 3780 383
<< metal1 >>
rect 0 724 4144 844
rect 201 703 247 724
rect 201 646 247 657
rect 498 703 544 724
rect 1424 703 1508 724
rect 498 646 544 657
rect 600 632 1124 678
rect 1424 657 1441 703
rect 1487 657 1508 703
rect 1896 703 1969 724
rect 1896 657 1909 703
rect 1955 657 1969 703
rect 2817 703 2863 724
rect 2431 666 2477 678
rect 600 600 646 632
rect 41 587 89 599
rect 221 587 646 600
rect 87 554 646 587
rect 693 574 739 585
rect 87 541 267 554
rect 41 530 89 541
rect 25 379 172 412
rect 25 333 113 379
rect 159 333 172 379
rect 25 320 172 333
rect 221 397 267 541
rect 349 453 361 499
rect 407 453 419 499
rect 221 378 281 397
rect 221 332 235 378
rect 221 321 281 332
rect 41 255 87 266
rect 221 255 267 321
rect 87 209 267 255
rect 361 255 407 453
rect 469 385 636 507
rect 469 339 590 385
rect 469 280 636 339
rect 682 468 693 506
rect 894 515 940 632
rect 682 457 739 468
rect 888 503 940 515
rect 360 209 361 234
rect 682 255 728 457
rect 888 439 940 451
rect 407 209 636 234
rect 41 198 87 209
rect 360 188 636 209
rect 682 198 728 209
rect 774 407 820 420
rect 590 152 636 188
rect 774 152 820 361
rect 894 371 940 439
rect 894 314 940 325
rect 986 569 1032 580
rect 986 273 1032 453
rect 1078 385 1124 632
rect 1182 622 1228 634
rect 1601 625 1647 636
rect 1228 579 1601 611
rect 1228 576 1647 579
rect 1182 565 1647 576
rect 1732 622 1778 633
rect 1778 576 1966 611
rect 1732 565 1966 576
rect 1078 326 1124 339
rect 1170 473 1857 519
rect 1170 273 1216 473
rect 1811 405 1857 473
rect 1367 391 1444 403
rect 986 255 1216 273
rect 1032 227 1216 255
rect 1263 347 1309 367
rect 1367 339 1378 391
rect 1430 358 1444 391
rect 1807 384 1871 405
rect 1920 403 1966 565
rect 2015 568 2382 608
rect 2015 562 2330 568
rect 1367 312 1387 339
rect 1433 312 1444 358
rect 1519 312 1530 358
rect 1576 312 1746 358
rect 1807 338 1818 384
rect 1864 338 1871 384
rect 1807 312 1871 338
rect 1917 391 1969 403
rect 1917 327 1969 339
rect 2015 384 2061 562
rect 2382 516 2385 567
rect 2015 325 2061 338
rect 2107 499 2159 510
rect 2107 453 2109 499
rect 2155 453 2159 499
rect 2107 391 2159 453
rect 2205 504 2257 516
rect 2330 514 2385 516
rect 2330 504 2382 514
rect 3186 703 3232 724
rect 2817 640 2863 653
rect 2909 630 3140 676
rect 3572 703 3618 724
rect 3186 642 3232 656
rect 2909 594 2955 630
rect 2477 548 2955 594
rect 3094 593 3140 630
rect 3278 632 3508 678
rect 3278 593 3324 632
rect 3001 572 3047 584
rect 2257 452 2385 458
rect 2205 406 2385 452
rect 2339 384 2385 406
rect 1263 263 1309 301
rect 1434 263 1446 266
rect 986 198 1032 209
rect 1263 217 1446 263
rect 1263 152 1309 217
rect 1434 214 1446 217
rect 1498 214 1510 266
rect 1700 259 1746 312
rect 1700 213 1947 259
rect 2107 255 2159 339
rect 201 127 247 138
rect 201 60 247 81
rect 498 127 544 138
rect 590 106 1309 152
rect 1901 152 1947 213
rect 2087 209 2098 255
rect 2144 209 2159 255
rect 2206 347 2258 360
rect 2206 301 2209 347
rect 2255 301 2258 347
rect 2339 325 2385 338
rect 2206 266 2258 301
rect 2431 255 2477 460
rect 2600 455 2611 501
rect 2657 455 2668 501
rect 2206 198 2258 214
rect 2304 209 2316 255
rect 2362 209 2477 255
rect 2524 403 2570 416
rect 2524 278 2570 357
rect 2524 266 2576 278
rect 2524 202 2576 214
rect 2622 265 2668 455
rect 2715 390 2945 502
rect 2715 338 2729 390
rect 2781 384 2945 390
rect 3094 547 3324 593
rect 3370 573 3416 585
rect 3001 384 3047 463
rect 2781 338 2888 384
rect 2934 338 2945 384
rect 2715 313 2945 338
rect 2994 333 3047 384
rect 3093 453 3370 493
rect 3093 447 3416 453
rect 3093 382 3139 447
rect 2994 265 3040 333
rect 3093 323 3139 336
rect 3191 347 3324 398
rect 2622 255 3040 265
rect 2622 209 2634 255
rect 2680 209 2809 255
rect 2855 209 3040 255
rect 3191 301 3267 347
rect 3313 301 3324 347
rect 3191 223 3324 301
rect 3370 315 3416 447
rect 3462 407 3508 632
rect 3572 429 3618 453
rect 3702 703 3748 724
rect 4022 703 4068 724
rect 3702 429 3748 453
rect 3843 667 3929 678
rect 3843 453 3862 667
rect 3908 453 3929 667
rect 3462 361 3473 407
rect 3519 361 3530 407
rect 3610 337 3624 383
rect 3780 337 3791 383
rect 3610 315 3656 337
rect 3370 269 3656 315
rect 3087 176 3324 223
rect 3554 255 3600 269
rect 3087 152 3134 176
rect 498 60 544 81
rect 1639 81 1651 127
rect 1697 81 1710 127
rect 1901 106 3134 152
rect 3554 141 3600 152
rect 3702 255 3748 278
rect 1639 60 1710 81
rect 3180 81 3195 127
rect 3241 81 3263 127
rect 3180 60 3263 81
rect 3843 255 3929 453
rect 4022 429 4068 453
rect 3843 117 3862 255
rect 3908 117 3929 255
rect 3843 106 3929 117
rect 4022 255 4068 277
rect 3702 60 3748 81
rect 4022 60 4068 81
rect 0 -60 4144 60
<< via1 >>
rect 888 451 940 503
rect 1378 358 1430 391
rect 1378 339 1387 358
rect 1387 339 1430 358
rect 1917 339 1969 391
rect 2330 516 2382 568
rect 2205 452 2257 504
rect 2107 339 2159 391
rect 1446 214 1498 266
rect 2206 214 2258 266
rect 2524 214 2576 266
rect 2729 338 2781 390
<< metal2 >>
rect 2327 568 2385 580
rect 2327 516 2330 568
rect 2382 516 2385 568
rect 2327 512 2385 516
rect 876 504 2270 506
rect 876 503 2205 504
rect 876 451 888 503
rect 940 452 2205 503
rect 2257 452 2270 504
rect 940 451 2270 452
rect 876 449 2270 451
rect 1366 391 2171 393
rect 1366 339 1378 391
rect 1430 339 1917 391
rect 1969 339 2107 391
rect 2159 339 2171 391
rect 1366 336 2171 339
rect 2329 392 2385 512
rect 2329 390 2793 392
rect 2329 338 2729 390
rect 2781 338 2793 390
rect 2329 336 2793 338
rect 1434 266 2589 268
rect 1434 214 1446 266
rect 1498 214 2206 266
rect 2258 214 2524 266
rect 2576 214 2589 266
rect 1434 212 2589 214
rect 1434 211 1502 212
<< labels >>
flabel metal1 s 0 724 4144 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 4144 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel metal1 25 320 172 412 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 3843 106 3929 678 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 s 3191 176 3324 398 0 FreeSans 416 0 0 0 RN
port 8 nsew
flabel metal1 s 2715 313 2945 502 0 FreeSans 416 0 0 0 SN
port 9 nsew
flabel metal1 s 469 280 636 507 0 FreeSans 416 0 0 0 D
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 4144 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 4160 354
string MASKHINTS_PPLUS -16 354 4160 830
<< end >>
